//Copyright (C)2014-2023 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//Tool Version: V1.9.9
//Part Number: GW2AR-LV18QN88C8/I7
//Device: GW2AR-18
//Device Version: C
//Created Time: Thu May 15 20:46:50 2025

module Gowin_SDPB (dout, clka, cea, reseta, clkb, ceb, resetb, oce, ada, din, adb);

output [1:0] dout;
input clka;
input cea;
input reseta;
input clkb;
input ceb;
input resetb;
input oce;
input [14:0] ada;
input [1:0] din;
input [14:0] adb;

wire [30:0] sdpb_inst_0_dout_w;
wire [0:0] sdpb_inst_0_dout;
wire [30:0] sdpb_inst_1_dout_w;
wire [0:0] sdpb_inst_1_dout;
wire [30:0] sdpb_inst_2_dout_w;
wire [1:1] sdpb_inst_2_dout;
wire [30:0] sdpb_inst_3_dout_w;
wire [1:1] sdpb_inst_3_dout;
wire dff_q_0;
wire gw_gnd;

assign gw_gnd = 1'b0;

SDPB sdpb_inst_0 (
    .DO({sdpb_inst_0_dout_w[30:0],sdpb_inst_0_dout[0]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({gw_gnd,gw_gnd,ada[14]}),
    .BLKSELB({gw_gnd,gw_gnd,adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[0]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_0.READ_MODE = 1'b0;
defparam sdpb_inst_0.BIT_WIDTH_0 = 1;
defparam sdpb_inst_0.BIT_WIDTH_1 = 1;
defparam sdpb_inst_0.BLK_SEL_0 = 3'b000;
defparam sdpb_inst_0.BLK_SEL_1 = 3'b000;
defparam sdpb_inst_0.RESET_MODE = "SYNC";
defparam sdpb_inst_0.INIT_RAM_00 = 256'h0000080800848902208100040000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_01 = 256'h0000804250100028082020802000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_02 = 256'h0000020428081060004004000000000BBF0FF790800000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_03 = 256'h000010200121890212048040000003BFFFFFFFFF980000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_04 = 256'h00000002284482008404000480003FFFFFFFFFFFFFD000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_05 = 256'h00004840010010640220210200003FFFFFFFFFFFFFFC00000000000000000000;
defparam sdpb_inst_0.INIT_RAM_06 = 256'h00001100801101051400044001007FFFFFFFFFFFFFFE00000000000000000000;
defparam sdpb_inst_0.INIT_RAM_07 = 256'h000000A2104488204061800000007FFFFFFFFFFFFFFC00000000000000000000;
defparam sdpb_inst_0.INIT_RAM_08 = 256'h00001202019129109811200000007FF7FFFFFFFFFFFE00000000000000000000;
defparam sdpb_inst_0.INIT_RAM_09 = 256'h00000020180800060100084412007FD9FFFFFFFFFFFC00000000000000000000;
defparam sdpb_inst_0.INIT_RAM_0A = 256'h00000000500091020080010000003F47FFFFFFFFFFFE00000000000000000000;
defparam sdpb_inst_0.INIT_RAM_0B = 256'h00004441021208900824801000023FF8FFFFFFFFFFFC00000000000000000000;
defparam sdpb_inst_0.INIT_RAM_0C = 256'h00001180229200209040018141507FF5FFFFFFFFFFFC00000000000000000000;
defparam sdpb_inst_0.INIT_RAM_0D = 256'h0000040A0800A50A0914582000007FCBFFFFFFFFFFFE00000000000000000000;
defparam sdpb_inst_0.INIT_RAM_0E = 256'h0000411490062482000A208408007FE5FFFFFFFFFFFE00000000000000000000;
defparam sdpb_inst_0.INIT_RAM_0F = 256'h00000000012000201440000110006FEBFFFFFFFFFFFF80000000000000000000;
defparam sdpb_inst_0.INIT_RAM_10 = 256'h0000186200009004A4240420800177EBFFFFFFFFFFFFFC000000000000000000;
defparam sdpb_inst_0.INIT_RAM_11 = 256'h0000000026660241000260040880FED7FFFFFFFFFFFFFC000000000000000000;
defparam sdpb_inst_0.INIT_RAM_12 = 256'h0000002052000A50895441002201FFEFFFFFFFFFFFFFFE000000000000000000;
defparam sdpb_inst_0.INIT_RAM_13 = 256'h0000440100429004100008820017FFFFFFFFFFFFFFFFFC000000000000000000;
defparam sdpb_inst_0.INIT_RAM_14 = 256'h00000808204A200904202110043FFFFFFFFFFFFFFFFFFE000000000000000000;
defparam sdpb_inst_0.INIT_RAM_15 = 256'h0000822102000A9020048082401FFFFFFFFFFFFFFFFFFC000000000000000000;
defparam sdpb_inst_0.INIT_RAM_16 = 256'h000004405A105009A6660004107FFFFFFFFFFFFFFFFFFC000000000000000000;
defparam sdpb_inst_0.INIT_RAM_17 = 256'h00001022004A052000001222040FFFFFFFFFFFFFFFFFFC000000000000000000;
defparam sdpb_inst_0.INIT_RAM_18 = 256'h00000022000A0A909000991484139FFFFFFFFFFFFFFF84000000000000000000;
defparam sdpb_inst_0.INIT_RAM_19 = 256'h000094809A4040090A660000101987FFFFFFFFFFFFFF8C000000000000000000;
defparam sdpb_inst_0.INIT_RAM_1A = 256'h000002090250559200000000005085FFFFFFFFFFFFFF8C000000000000000000;
defparam sdpb_inst_0.INIT_RAM_1B = 256'h00000820400A000094422819411103FEFFFFF0FFFFFF04000000000000000000;
defparam sdpb_inst_0.INIT_RAM_1C = 256'h0000000490000000054A91901012807FFFFFF9FFFFEF04000000000000000000;
defparam sdpb_inst_0.INIT_RAM_1D = 256'h0000A2200296A56A9000000088927B9FFFFFF8FFFFDF8C000000000000000000;
defparam sdpb_inst_0.INIT_RAM_1E = 256'h000006A619801002201008000C91FFFFFFFFF9FFFFFFFC000000000000000000;
defparam sdpb_inst_0.INIT_RAM_1F = 256'h0000400080150950054A919E2957BFFFFFFFF1FFFFFFFC000000000000000000;
defparam sdpb_inst_0.INIT_RAM_20 = 256'h00002000004128180A2007AFD2FCBFFFFFFFFFFFFFFFFC000000000000000000;
defparam sdpb_inst_0.INIT_RAM_21 = 256'h0000059696284181400DD11FFE6B7FFFFFFFF1FFFFFF07A00000000000000000;
defparam sdpb_inst_0.INIT_RAM_22 = 256'h0000540000050A5990DFFFDFFF10FFFAFFFFE3FFFFF18A08F800000000000000;
defparam sdpb_inst_0.INIT_RAM_23 = 256'h0000009295A050000BFF8DFFFF8AFFFF114FF5FFBFBF97D74387900000000000;
defparam sdpb_inst_0.INIT_RAM_24 = 256'h000020011051204411A0FAFFFFD7FFFFABFEE3F0BFFFBFF7EFFFEA3800000000;
defparam sdpb_inst_0.INIT_RAM_25 = 256'h0000052481084522891279FFFFFEFFFFFFFFE17F47FFFFFFFDAA007E00000000;
defparam sdpb_inst_0.INIT_RAM_26 = 256'h000064805A450800910E7FFFFFCFFFFFFBCFE042EFFFFFFFFB7FFBEC00000000;
defparam sdpb_inst_0.INIT_RAM_27 = 256'h00000025002051AA082C3FFFFE7AFFFF047FF93FFBFFFFFFFFFFD7E000000000;
defparam sdpb_inst_0.INIT_RAM_28 = 256'h00000100004A04AA14013FFFFAF2FFFFC977F0FFFFFFDFFFEFA2BFD000000000;
defparam sdpb_inst_0.INIT_RAM_29 = 256'h00006455AA10A10042A4FBDFF9AFFFF5FEDFF7FEFF7FE860305F65EC00000000;
defparam sdpb_inst_0.INIT_RAM_2A = 256'h0000004811021A2210017FFFF9D2FFF6770BFFFFFFDF7FAB6FFDC8F800000000;
defparam sdpb_inst_0.INIT_RAM_2B = 256'h0000451089AC804444957FBFFEBCFFF67D3E1B5FFFFFDBF6502137DC00000000;
defparam sdpb_inst_0.INIT_RAM_2C = 256'h00005A13426480150A20FFF7FDFAFFFB6A100A138042FFFAAD9BC09C00000000;
defparam sdpb_inst_0.INIT_RAM_2D = 256'h0000008424021D80504D7EF3FEA5FFFFFFFFDCCC8100BA282BC0009800000000;
defparam sdpb_inst_0.INIT_RAM_2E = 256'h0000A0500168805441FEFFF7FDA4FFFFFFFFFFFFFF9A16FAD10102DC00000000;
defparam sdpb_inst_0.INIT_RAM_2F = 256'h00000605A402290313FF7FC7F829FFFFFFFFFFFFFF9EFFC40000009800000000;
defparam sdpb_inst_0.INIT_RAM_30 = 256'h000041042104A0503FFFFFFFFF99FFFFFFFFFFFFFFBA04008842029800000000;
defparam sdpb_inst_0.INIT_RAM_31 = 256'h000028A188A1850BFFFFFFFFFFFFFFFFFFFFFFFFFFDC6048000000FC01000400;
defparam sdpb_inst_0.INIT_RAM_32 = 256'h00000512012A511FFFFFFFFFFFFFFFFFFFFFFFFFFF9F40822120009C00810000;
defparam sdpb_inst_0.INIT_RAM_33 = 256'h0000A08854800A7FFFFFFFFFFFFFFFFFFFFFFFFFFF9FFFA0000820D840000000;
defparam sdpb_inst_0.INIT_RAM_34 = 256'h000001081C80044217FFFFFFFFFFFFFFFFFFFFFFFFBB4BCFFFB0009804000000;
defparam sdpb_inst_0.INIT_RAM_35 = 256'h000058A24215A40087FFFFFFFFFFFFFFFFFFFFFFFFDEFEA65FFFDF3C00800104;
defparam sdpb_inst_0.INIT_RAM_36 = 256'h000081218848125827FFFFFFFFFFFFFFFFFFFFFFFFDEDF07F5E77FB8F4008040;
defparam sdpb_inst_0.INIT_RAM_37 = 256'h00001484212993E103EFFFFFFFFFFFFFFFFFFFFFFF9DE95D8BD0621B8FCE2000;
defparam sdpb_inst_0.INIT_RAM_38 = 256'h0000A503C2C047E483FFFFFFFFFFFFFFFFFFFFFFFFDF0A5FA5D7D4BCAE1C2004;
defparam sdpb_inst_0.INIT_RAM_39 = 256'h00000054242A3FE01DFFFFFFFFFFFFFFFFFFFFFFFF9F8FA26A17FFF2AEF80210;
defparam sdpb_inst_0.INIT_RAM_3A = 256'h0000248181827FE001FFFFFFFFFFFFFFFFFFFFFFFFDFFFF356FFFFFFFFF20082;
defparam sdpb_inst_0.INIT_RAM_3B = 256'h0000A21424283DE805FFFEFFFFFFFFFFFFFFFFFFFF9FFF3524FFFBFEBF824800;
defparam sdpb_inst_0.INIT_RAM_3C = 256'h000011042422612695FFFFFFFFFFFBFFFFFFFFFFFF9F95AB57FF128FFF4C1000;
defparam sdpb_inst_0.INIT_RAM_3D = 256'h000088624244046607FFFFFFFFFFFFFFFFFFFFF7FF98B971FFFF77307A228218;
defparam sdpb_inst_0.INIT_RAM_3E = 256'h000055000000087003FFFFFFFFFFFFFFFFFFFFF7FE3C62BFFFFFC360AAA00000;
defparam sdpb_inst_0.INIT_RAM_3F = 256'h000000AA5A55936727FFFFFFFFFFF3FFFFFFFFFFFF3EDFFFFFFF863DD2042481;

SDPB sdpb_inst_1 (
    .DO({sdpb_inst_1_dout_w[30:0],sdpb_inst_1_dout[0]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({gw_gnd,gw_gnd,ada[14]}),
    .BLKSELB({gw_gnd,gw_gnd,adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[0]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_1.READ_MODE = 1'b0;
defparam sdpb_inst_1.BIT_WIDTH_0 = 1;
defparam sdpb_inst_1.BIT_WIDTH_1 = 1;
defparam sdpb_inst_1.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_1.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_1.RESET_MODE = "SYNC";
defparam sdpb_inst_1.INIT_RAM_00 = 256'h00000A500950457DA7FFFFFFFFFFFFFFFFFFFFEBFF3FFFFFFFD9835BBC080182;
defparam sdpb_inst_1.INIT_RAM_01 = 256'h00005004A0051DF01FFCFFFFFFFFFBFFFFD7FFFDF87FFFFFFFBF82EF0C214800;
defparam sdpb_inst_1.INIT_RAM_02 = 256'h0000400910084DF80FF87FFFFFFFFFFFFF5639A7FE7FFFED9F2A93BE55402014;
defparam sdpb_inst_1.INIT_RAM_03 = 256'h00000A5005501B612FF7FFDFFFC37FFFFFFFFFD9ADFFFFBBFE1F83EA43208000;
defparam sdpb_inst_1.INIT_RAM_04 = 256'h00000249844916E41DFBFFFFFFFFFFFFFFFFCCED15FBFD7BBF0EC3D9AB100081;
defparam sdpb_inst_1.INIT_RAM_05 = 256'h00004000100046F07DFBFFFFFFCBFFFFBEA7FFFEEAFFFFFDFE9D497071021124;
defparam sdpb_inst_1.INIT_RAM_06 = 256'h00002820002011E1FFDFFFFFFFFFFFFD38ED1E67FF1FF647F98093E045888401;
defparam sdpb_inst_1.INIT_RAM_07 = 256'h00008084488436E8FFF3FF2FFF5BFFFF8029E27340197FF9FC1FA3045AC00080;
defparam sdpb_inst_1.INIT_RAM_08 = 256'h00000040102039E9FFFFFFEFFFBCFFFFFFFCF48EB4304FEFFB742F8073C60440;
defparam sdpb_inst_1.INIT_RAM_09 = 256'h0000080A800263DFFFCFFE1FFC97FFFD7BFEFEDF75A45FD565FC620BDE400000;
defparam sdpb_inst_1.INIT_RAM_0A = 256'h00004010020821E7FFFFFD3FFFBBFFDF7FFFFFFFFE1FDF7DE67C2400BFC02000;
defparam sdpb_inst_1.INIT_RAM_0B = 256'h0000020000200563FFFFF01FF301FFA9CBFFEDFFFFFFEDDBD5BCDE01DCE00808;
defparam sdpb_inst_1.INIT_RAM_0C = 256'h00000001000095CFFFFFF87FFB23FF3BBFFFB796BA55FFEFF98C6C41F1600040;
defparam sdpb_inst_1.INIT_RAM_0D = 256'h00000000000001EFF6FFFA7FF10BFF3093FDC7F96BFFBFB5FFAD2C07E4200000;
defparam sdpb_inst_1.INIT_RAM_0E = 256'h00000000000023FFF0FFF3FFCC4FFC2F07FC7BCEE685BF87FA97780AFA600000;
defparam sdpb_inst_1.INIT_RAM_0F = 256'h0000000000001DDFF07FD0FFD01FFF2A5FFA1A44556A1ED7FF4B183FE0200000;
defparam sdpb_inst_1.INIT_RAM_10 = 256'h00000000000037FFE1FF93FF9BBFFB754FFA98A01915BF9FFF87FE3761200000;
defparam sdpb_inst_1.INIT_RAM_11 = 256'h0000000000003BFF83FFDFFF283FF43A97F9C2F80F3B1E77F7FBFFFF60200000;
defparam sdpb_inst_1.INIT_RAM_12 = 256'h00000000000033FF83FFCFFF62BFE1B56FFED5DEFC338C8FFFF9FFFC66380000;
defparam sdpb_inst_1.INIT_RAM_13 = 256'h00000000000007FF03FFDFFF9EFFF43C2FFEAB765C354D3F9DCFEFFEE02C0000;
defparam sdpb_inst_1.INIT_RAM_14 = 256'h0000000000001FFE07FFDFFF3DFFD6AF87F9278954043D6FDDA9BFFFEFB80000;
defparam sdpb_inst_1.INIT_RAM_15 = 256'h00000000000003FE0FFFDFFFFEFF2BDAB9FF207AA6D74E177FFDCBFFEF200000;
defparam sdpb_inst_1.INIT_RAM_16 = 256'h0000000000001FFC0FF39FFFFFEF14FFFF55F7D4DA25BD1FCFFFABFEBE800000;
defparam sdpb_inst_1.INIT_RAM_17 = 256'h0000000000000FFC3FF39FFEF5FFFF1071F4AA69E4931EEFFF7BBDFC5E300000;
defparam sdpb_inst_1.INIT_RAM_18 = 256'h0000000000001FF07FF7FFFFFFFFFFFFFFFFFFF52043BF6FBFEDFFFF9A400000;
defparam sdpb_inst_1.INIT_RAM_19 = 256'h0000000000000FF07FF2FFFFFFFEEBFFFFFBB7855511DC5FDFE3FFFFC0400000;
defparam sdpb_inst_1.INIT_RAM_1A = 256'h0000000000003FF87FEDFFFFFFFFFEF6FFFF900AFFFF3E57BF539DFF81000000;
defparam sdpb_inst_1.INIT_RAM_1B = 256'h0000000000007FFCFF40FFFBFFFFFFBFFFFFFFFD0FFFBF9FEDEF8FFC89C00000;
defparam sdpb_inst_1.INIT_RAM_1C = 256'h000000000000FF7FFFC7FFBDFFFFFFFD6A1BDB09BEFFBEAFFFAFA7FD54800000;
defparam sdpb_inst_1.INIT_RAM_1D = 256'h0000000000007F413F6FFEFF3FFFEFC853DFEFFFE7FFBFAFA957DFFDA5000000;
defparam sdpb_inst_1.INIT_RAM_1E = 256'h000000000000BF85801FFEE77FFA2FFF79EFFFFFFFFFBB2FFDA7E3C449800000;
defparam sdpb_inst_1.INIT_RAM_1F = 256'h0000000000003FFB803F9FB3FFFFC2FFAFFFFFDFDDFFFABED74FEBB0D7000000;
defparam sdpb_inst_1.INIT_RAM_20 = 256'h0000000000001FFFF81FFFC0FF2FFFFC6F0BFFEFBFFC3BDF7ECFE1D0D5000000;
defparam sdpb_inst_1.INIT_RAM_21 = 256'h0000000000001FFFF03FF780EF009FBC79EC3C4FFFFFD337697D703E2A000000;
defparam sdpb_inst_1.INIT_RAM_22 = 256'h0000000000000FFFFE3FE403FE000005F00786F80200BE5FBA7C284F76000000;
defparam sdpb_inst_1.INIT_RAM_23 = 256'h0000000000000FFFFEBFFC039E000000002F8028800577EDF7F81003F8000000;
defparam sdpb_inst_1.INIT_RAM_24 = 256'h0000000000000FFFEFFFC00FFC00000000000057F2941F3FDFD80006E8000000;
defparam sdpb_inst_1.INIT_RAM_25 = 256'h0000000000000FFF9FFFC00770000000000000000001948BA908300998000000;
defparam sdpb_inst_1.INIT_RAM_26 = 256'h0000000000000FFF001FE01EF0000000000000000000003FFB08230BF0000000;
defparam sdpb_inst_1.INIT_RAM_27 = 256'h0000000000001FFE001FE01EE00000000000000000000005FE08031D40000000;
defparam sdpb_inst_1.INIT_RAM_28 = 256'h0000000000001FFE001FC07DE0000000000000000000000BF808012FC0000000;
defparam sdpb_inst_1.INIT_RAM_29 = 256'h0000000000001FFC003FC07BC00000000000000000000008F808096980000000;
defparam sdpb_inst_1.INIT_RAM_2A = 256'h0000000000001FFC001FC0F7800000000000000000000006FC4821DF00000000;
defparam sdpb_inst_1.INIT_RAM_2B = 256'h0000000000001FF0001FC0F78000000000000000000000023E0807F600000000;
defparam sdpb_inst_1.INIT_RAM_2C = 256'h0000000000003FE0003FC1EF0000000000000000000000002E0411FC00000000;
defparam sdpb_inst_1.INIT_RAM_2D = 256'h0000000000003FF0001FE1FF0000000000000000000000005FC87FF000000000;
defparam sdpb_inst_1.INIT_RAM_2E = 256'h0000000000007FE0001FC3DC0000000000000000000000001FFFFFC000000000;
defparam sdpb_inst_1.INIT_RAM_2F = 256'h0000000000007FC0001FC7B800000000000000000000000007FFFF0000000000;
defparam sdpb_inst_1.INIT_RAM_30 = 256'h000000000000FFE0003FCF7000000000000000000000000000DFD00000000000;
defparam sdpb_inst_1.INIT_RAM_31 = 256'h000000000000FFE0003FDEF00000000000000000000000000000000000000000;
defparam sdpb_inst_1.INIT_RAM_32 = 256'h000000000001FFC0003FFEF00000000000000000000000000000000000000000;
defparam sdpb_inst_1.INIT_RAM_33 = 256'h000000000001FFE0001FFFE00000000000000000000000000000000000000000;
defparam sdpb_inst_1.INIT_RAM_34 = 256'h000000000003FFFD8C7FFFC00000000000000000000000000000000000000000;
defparam sdpb_inst_1.INIT_RAM_35 = 256'h000000000003FFFFDFFFFF800000000000000000000000000000000000000000;
defparam sdpb_inst_1.INIT_RAM_36 = 256'h000000000003FFFFFFFFFF800000000000000000000000000000000000000000;
defparam sdpb_inst_1.INIT_RAM_37 = 256'h000000000003FFFFDFFFFF000000000000000000000000000000000000000000;
defparam sdpb_inst_1.INIT_RAM_38 = 256'h0000000000B3FFE01FFFFF000000000000000000000000000000000000000000;
defparam sdpb_inst_1.INIT_RAM_39 = 256'h0000000006FFFC009DFFFC000000000000000000000000000000000000000000;
defparam sdpb_inst_1.INIT_RAM_3A = 256'h00000006FFFF573FFFC754000000000000000000000000000000000000000000;
defparam sdpb_inst_1.INIT_RAM_3B = 256'h00000003FFFFFFFFFE0000000000000000000000000000000000000000000000;
defparam sdpb_inst_1.INIT_RAM_3C = 256'h000000006E3FFFEC000000000000000000000000000000000000000000000000;
defparam sdpb_inst_1.INIT_RAM_3D = 256'h00000000000A9A80000000000000000000000000000000000000000000000000;

SDPB sdpb_inst_2 (
    .DO({sdpb_inst_2_dout_w[30:0],sdpb_inst_2_dout[1]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({gw_gnd,gw_gnd,ada[14]}),
    .BLKSELB({gw_gnd,gw_gnd,adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[1]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_2.READ_MODE = 1'b0;
defparam sdpb_inst_2.BIT_WIDTH_0 = 1;
defparam sdpb_inst_2.BIT_WIDTH_1 = 1;
defparam sdpb_inst_2.BLK_SEL_0 = 3'b000;
defparam sdpb_inst_2.BLK_SEL_1 = 3'b000;
defparam sdpb_inst_2.RESET_MODE = "SYNC";
defparam sdpb_inst_2.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_2.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_2.INIT_RAM_02 = 256'h0000000000000000000000000000000000F00800000000000000000000000000;
defparam sdpb_inst_2.INIT_RAM_03 = 256'h0000000000000000000000000000007FFFFFFFFFE00000000000000000000000;
defparam sdpb_inst_2.INIT_RAM_04 = 256'h00000000000000000000000000001FFFFFFFFFFFFFE000000000000000000000;
defparam sdpb_inst_2.INIT_RAM_05 = 256'h00000000000000000000000000003FFFFFFFFFFFFFF800000000000000000000;
defparam sdpb_inst_2.INIT_RAM_06 = 256'h00000000000000000000000000003FFFFFFFFFFFFFFC00000000000000000000;
defparam sdpb_inst_2.INIT_RAM_07 = 256'h00000000000000000000000000003FFFFFFFFFFFFFFE00000000000000000000;
defparam sdpb_inst_2.INIT_RAM_08 = 256'h00000000000000000000000000003FFFFFFFFFFFFFFC00000000000000000000;
defparam sdpb_inst_2.INIT_RAM_09 = 256'h00000000000000000000000000003FFFFFFFFFFFFFFC00000000000000000000;
defparam sdpb_inst_2.INIT_RAM_0A = 256'h00000000000000000000000000007FFFFFFFFFFFFFFC00000000000000000000;
defparam sdpb_inst_2.INIT_RAM_0B = 256'h00000000000000000000000000007F7FFFFFFFFFFFFE00000000000000000000;
defparam sdpb_inst_2.INIT_RAM_0C = 256'h00000000000000000000000000007FFFFFFFFFFFFFFC00000000000000000000;
defparam sdpb_inst_2.INIT_RAM_0D = 256'h00000000000000000000000000007FFFFFFFFFFFFFFC00000000000000000000;
defparam sdpb_inst_2.INIT_RAM_0E = 256'h00000000000000000000000000007FFFFFFFFFFFFFFC00000000000000000000;
defparam sdpb_inst_2.INIT_RAM_0F = 256'h00000000000000000000000000007FFFFFFFFFFFFFFF00000000000000000000;
defparam sdpb_inst_2.INIT_RAM_10 = 256'h00000000000000000000000000007FFFFFFFFFFFFFFFF8000000000000000000;
defparam sdpb_inst_2.INIT_RAM_11 = 256'h00000000000000000000000000007FFFFFFFFFFFFFFFFC000000000000000000;
defparam sdpb_inst_2.INIT_RAM_12 = 256'h0000000000000000000000000000FFFFFFFFFFFFFFFFFC000000000000000000;
defparam sdpb_inst_2.INIT_RAM_13 = 256'h000000000000000000000000000FFFFFFFFFFFFFFFFFFE000000000000000000;
defparam sdpb_inst_2.INIT_RAM_14 = 256'h000000000000000000000000001FFFFFFFFFFFFFFFFFFC000000000000000000;
defparam sdpb_inst_2.INIT_RAM_15 = 256'h000000000000000000000000001FFFFFFFFFFFFFFFFFFC000000000000000000;
defparam sdpb_inst_2.INIT_RAM_16 = 256'h000000000000000000000000001FFFFFFFFFFFFFFFFFF8000000000000000000;
defparam sdpb_inst_2.INIT_RAM_17 = 256'h000000000000000000000000001FFFFFFFFFFFFFFFFFF8000000000000000000;
defparam sdpb_inst_2.INIT_RAM_18 = 256'h000000000000000000000000000F03FFFFFFFFFFFFFFF8000000000000000000;
defparam sdpb_inst_2.INIT_RAM_19 = 256'h000000000000000000000000000F03FFFFFFFFFFFFFFF8000000000000000000;
defparam sdpb_inst_2.INIT_RAM_1A = 256'h000000000000000000000000000F03FFFFFFFFFFFFFFF8000000000000000000;
defparam sdpb_inst_2.INIT_RAM_1B = 256'h000000000000000000000000000F00FFFFFFFFFFFFFFF8000000000000000000;
defparam sdpb_inst_2.INIT_RAM_1C = 256'h000000000000000000000000000F000FFFFFF7FFFFFFF8000000000000000000;
defparam sdpb_inst_2.INIT_RAM_1D = 256'h000000000000000000000000000F00FFFFFFF7FFFFFFF8000000000000000000;
defparam sdpb_inst_2.INIT_RAM_1E = 256'h000000000000000000000000026FFFFFFFFFC7FFFFFFFC000000000000000000;
defparam sdpb_inst_2.INIT_RAM_1F = 256'h000000000000000000000001FE007FFFFFFFFFFFFFFFF8000000000000000000;
defparam sdpb_inst_2.INIT_RAM_20 = 256'h00000000000000000000007FFF007FFFFFFFF1FFFFFFF8000000000000000000;
defparam sdpb_inst_2.INIT_RAM_21 = 256'h000000000000000000003EFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000;
defparam sdpb_inst_2.INIT_RAM_22 = 256'h0000000000000000003FFFFFFFFFFFFDFFFFFDFFFFFF7DF70000000000000000;
defparam sdpb_inst_2.INIT_RAM_23 = 256'h000000000000000000FFFFFFFFFFFFFFEFFFFFFFFFFF7FFFFFF8000000000000;
defparam sdpb_inst_2.INIT_RAM_24 = 256'h000000000000000000DFFFFFF83FFFFFFFFFDFFFFFFFFFFFFFFFFFC000000000;
defparam sdpb_inst_2.INIT_RAM_25 = 256'h000000000000000000ED87FFF807FFFFFFFFFFFFFFFFFFFFFFFDFFFE00000000;
defparam sdpb_inst_2.INIT_RAM_26 = 256'h000000000000000000F180FFFFE7FFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000;
defparam sdpb_inst_2.INIT_RAM_27 = 256'h00000000000000000001E0FFFFE7FFFFFFFFE7FFFFFFFFFFFFFFFFFE00000000;
defparam sdpb_inst_2.INIT_RAM_28 = 256'h00000000000000000000F3FFFFEFFFFFFFFFEFFFFFFFFFFFFFFFFFFE00000000;
defparam sdpb_inst_2.INIT_RAM_29 = 256'h0000000000000000000173FFFFC7FFFBFFFFFFFFFFFFFFFFFFFFFFF800000000;
defparam sdpb_inst_2.INIT_RAM_2A = 256'h00000000000000000000F3FFFE0FFFF988FFFFFFFFFFFFFFFFFFFFF800000000;
defparam sdpb_inst_2.INIT_RAM_2B = 256'h00000000000000000000FFFFFFFFFFF982C1FFFFFFFFFFFFFFFFF83800000000;
defparam sdpb_inst_2.INIT_RAM_2C = 256'h000000000000000000017FFFFFFFFFF7FFFFFFECFFFFFFFFF7FC007800000000;
defparam sdpb_inst_2.INIT_RAM_2D = 256'h00000000000000000000FFF7FFFFFFF7FFFFFFFFFFFF6FFFFC00007800000000;
defparam sdpb_inst_2.INIT_RAM_2E = 256'h0000000000000000003F7FE7FFFFFFFFFFFFFFFFFFFFFFFF0000003800000000;
defparam sdpb_inst_2.INIT_RAM_2F = 256'h000000000000000007FFFFE7FFFFFFFFFFFFFFFFFFFC00000000007800000000;
defparam sdpb_inst_2.INIT_RAM_30 = 256'h00000000000000001FFFFFC7FFEFFFFFFFFFFFFFFFDC00000000007800000000;
defparam sdpb_inst_2.INIT_RAM_31 = 256'h00000000000000007FFFFFF7FFFFFFFFFFFFFFFFFFF800000000003800000000;
defparam sdpb_inst_2.INIT_RAM_32 = 256'h00000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFCFF000000007800000000;
defparam sdpb_inst_2.INIT_RAM_33 = 256'h00000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000003800000000;
defparam sdpb_inst_2.INIT_RAM_34 = 256'h00000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFDCFFF00000007800000000;
defparam sdpb_inst_2.INIT_RAM_35 = 256'h00000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFC7FFFFFFFE0F800000000;
defparam sdpb_inst_2.INIT_RAM_36 = 256'h00000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00FFFFFFFFFF00000000;
defparam sdpb_inst_2.INIT_RAM_37 = 256'h00000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0007FFFFFDFF7FF00000;
defparam sdpb_inst_2.INIT_RAM_38 = 256'h0000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFCC007FFFFFF7FFFFE0000;
defparam sdpb_inst_2.INIT_RAM_39 = 256'h0000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00FFFFFFFFFFFFE0000;
defparam sdpb_inst_2.INIT_RAM_3A = 256'h0000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0FFFFFFFFFFFFC0000;
defparam sdpb_inst_2.INIT_RAM_3B = 256'h00000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDEFFFFFFFFFFFFC0000;
defparam sdpb_inst_2.INIT_RAM_3C = 256'h00000000000007FBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFFFFF00000;
defparam sdpb_inst_2.INIT_RAM_3D = 256'h00000000000007DDFFFFFFFFFFFFF3FFFFFFFFFFFFFFF7BFFFFFEBFFFFC00000;
defparam sdpb_inst_2.INIT_RAM_3E = 256'h00000000000007DFFFFFFFFFFFFFF3FFFFFFFFFFFFFFFFFFFFFFFFBF7D000000;
defparam sdpb_inst_2.INIT_RAM_3F = 256'h00000000000007FDFFFFFFFFFFFFFFFFFFFFFFF7FFFDFFFFFFFFFBFFFC000000;

SDPB sdpb_inst_3 (
    .DO({sdpb_inst_3_dout_w[30:0],sdpb_inst_3_dout[1]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({gw_gnd,gw_gnd,ada[14]}),
    .BLKSELB({gw_gnd,gw_gnd,adb[14]}),
    .ADA(ada[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[1]}),
    .ADB(adb[13:0])
);

defparam sdpb_inst_3.READ_MODE = 1'b0;
defparam sdpb_inst_3.BIT_WIDTH_0 = 1;
defparam sdpb_inst_3.BIT_WIDTH_1 = 1;
defparam sdpb_inst_3.BLK_SEL_0 = 3'b001;
defparam sdpb_inst_3.BLK_SEL_1 = 3'b001;
defparam sdpb_inst_3.RESET_MODE = "SYNC";
defparam sdpb_inst_3.INIT_RAM_00 = 256'h00000000000007F80FFFFFFFFFFFFFFFFFFFFFF7FFFFFFFFFFFFFFFFE8000000;
defparam sdpb_inst_3.INIT_RAM_01 = 256'h00000000000007F807FF3FFFFFFFFFFFFFFFFFE7FFBFFFFFFFDFFFFFFC000000;
defparam sdpb_inst_3.INIT_RAM_02 = 256'h0000000000000FF00FFFFFFFFFFFFFFFFFFFFFFFFFBFFFFFFFDFEFFFBE000000;
defparam sdpb_inst_3.INIT_RAM_03 = 256'h0000000000000FF01FFBFFFFFFFFFFFFFFFFFFFFFFBFFFFFFFFFFFFDFE000000;
defparam sdpb_inst_3.INIT_RAM_04 = 256'h0000000000000BF03FFFFFFFFF803FFFFFEFFFFFFEBFFFFFFFFFFFF0FF000000;
defparam sdpb_inst_3.INIT_RAM_05 = 256'h0000000000001FE03FFFFFFFFFBC3FFFF95FFFFFFF3FFFFFFF77F7E1FF800000;
defparam sdpb_inst_3.INIT_RAM_06 = 256'h0000000000001FE07FFBFFFFFFFFFFFAC712FBBFFFFFFFFFFF7FEFC1FF800000;
defparam sdpb_inst_3.INIT_RAM_07 = 256'h0000000000001FF0FFFFFFFFFFFFFFFFFFD61F8DBFF7FFFFFFFC3F81FF800000;
defparam sdpb_inst_3.INIT_RAM_08 = 256'h00000000000017FFFFFFFFFFFFFFFFFFFFFF1F754BDFFFFFFF9C3F01FFC00000;
defparam sdpb_inst_3.INIT_RAM_09 = 256'h0000000000001FFFFFFFFFFFFFFFFFFFFFFC3FFFFFFFFFFFFFFC3E007FC00000;
defparam sdpb_inst_3.INIT_RAM_0A = 256'h0000000000001FCFFFFFFACFFFFFFFFFFFFFFFFFFFE03C3FFFFC7E01FFC00000;
defparam sdpb_inst_3.INIT_RAM_0B = 256'h0000000000003FC7FFFFFFFFFCFFFFFFFFFFFFFFFFFFDE3FFFFC7C01FFC00000;
defparam sdpb_inst_3.INIT_RAM_0C = 256'h0000000000003FC7FFFFFFFFF4DFFFFFFFFFFFFFFFFFDFFFFFFCFC03FFC00000;
defparam sdpb_inst_3.INIT_RAM_0D = 256'h0000000000003FCFF9FFFFFFFFFFFFFF6FFFFFFFFFFFDFFFFFFCF807FFE00000;
defparam sdpb_inst_3.INIT_RAM_0E = 256'h0000000000003FCFF07FDFFFFFFFFFF0FFFFBFFFFFFFDFFFFFFEF80FFFE00000;
defparam sdpb_inst_3.INIT_RAM_0F = 256'h00000000000037FFE0FFFFFFFFFFFFF5BFFFE7BBBFFFFFFFFFFFF01FFFE00000;
defparam sdpb_inst_3.INIT_RAM_10 = 256'h0000000000001FFFC0FFFFFFFFFFFFFFFFFD67FFEFFFDFFFFFFFF03FFEE00000;
defparam sdpb_inst_3.INIT_RAM_11 = 256'h0000000000001FFFC1FFBFFFFFFFFFFFFFFE3F07F0C4FFAFFFFFFFFEFFE00000;
defparam sdpb_inst_3.INIT_RAM_12 = 256'h0000000000001FFF83FFBFFFFFFFFFFFFFFFFF2103CC7FFFFFFFFFFFF9E00000;
defparam sdpb_inst_3.INIT_RAM_13 = 256'h0000000000001FFF07FFBFFFE1FFFFDBFFFFFFFFFFFFFFFFE2FFFFFF7FFC0000;
defparam sdpb_inst_3.INIT_RAM_14 = 256'h0000000000001FFF0FFFBFFFE2FFFFFFFFFFFFFFFFFFDFBFE2FFFFFFF07C0000;
defparam sdpb_inst_3.INIT_RAM_15 = 256'h0000000000001FFE0FFBBFFFFFFFFFFFFFFEDFFFFFFDFFFFFFFFFFFFF0FC0000;
defparam sdpb_inst_3.INIT_RAM_16 = 256'h0000000000000FFC1FFFFFFFFFFFFFFFFFBFFFAB7FFFDFFFFFFFFFFFFD7C0000;
defparam sdpb_inst_3.INIT_RAM_17 = 256'h0000000000000FF81FEFFFFFFFFFFFFFFFFFFDFF9FFEFFBFFFFFFFFFFFE00000;
defparam sdpb_inst_3.INIT_RAM_18 = 256'h0000000000000FF83FFBFFFFFFFFFFFFFFFFFFFFFFFFDFBFFFFFFFFFFFC00000;
defparam sdpb_inst_3.INIT_RAM_19 = 256'h0000000000001FF87FFFFFFFFFFFFFFFFFFFFFFFFFFE7FFFFFFFFFFFFFC00000;
defparam sdpb_inst_3.INIT_RAM_1A = 256'h0000000000001FF8FF97FFFFFFFFFFFFFFFFFFF7FFFFDFFFFFFFFFFFFFC00000;
defparam sdpb_inst_3.INIT_RAM_1B = 256'h0000000000003FFCFFBFFFFFFFFFFFFFFFFFFFFFFFFFDFFFFFFFFFFFFF800000;
defparam sdpb_inst_3.INIT_RAM_1C = 256'h000000000000FFFDFFBFFF03FFFFFFFFFFFFFFFFFFFFDFFFFFFFFFFFFF800000;
defparam sdpb_inst_3.INIT_RAM_1D = 256'h000000000000FFBFFFFFFF00FFFFFFFFFFFFFFFFFFFFDFFFFFFFFFFE7F800000;
defparam sdpb_inst_3.INIT_RAM_1E = 256'h0000000000007FFA7FFFFF08FFC1FFFFFFFFFFFFFFFFDFFFFFFFFFF8FF000000;
defparam sdpb_inst_3.INIT_RAM_1F = 256'h0000000000003FFFFFDFFFE0FFC03D03FFFFFFFFFFFFDFFFFFFFFFE0FF000000;
defparam sdpb_inst_3.INIT_RAM_20 = 256'h0000000000001FFFF3FFFF80FF98000390FFFFFFFFFFDFFFFFFFFFE1FE000000;
defparam sdpb_inst_3.INIT_RAM_21 = 256'h0000000000001FFFF3FFFF01FF0000438613FFFFFFFFFFFFFFFFEFF9FE000000;
defparam sdpb_inst_3.INIT_RAM_22 = 256'h0000000000001FFFF1FFFE01DE0000000FF87F07FDFFFFFFFFF8173FFC000000;
defparam sdpb_inst_3.INIT_RAM_23 = 256'h0000000000001FFFFFFFF803FC00000000007FFF7FFADFFFFFE81F0FFC000000;
defparam sdpb_inst_3.INIT_RAM_24 = 256'h0000000000001FFBFFFFE007B8000000000000000FFFFFFF8FE81F07F8000000;
defparam sdpb_inst_3.INIT_RAM_25 = 256'h0000000000001FF787FFC00FF8000000000000000000003FDFF80F0FF0000000;
defparam sdpb_inst_3.INIT_RAM_26 = 256'h0000000000001FFF001FC00FF0000000000000000000001FFEF81D1FF0000000;
defparam sdpb_inst_3.INIT_RAM_27 = 256'h0000000000001FEF001FC01FF0000000000000000000001FFCF81D3FE0000000;
defparam sdpb_inst_3.INIT_RAM_28 = 256'h0000000000001FFE001FC03FC0000000000000000000000FF8F81F7FC0000000;
defparam sdpb_inst_3.INIT_RAM_29 = 256'h0000000000001FFC001FC03FC00000000000000000000007F0F817FF80000000;
defparam sdpb_inst_3.INIT_RAM_2A = 256'h0000000000001FF8001FC07F800000000000000000000003F8B81FFF00000000;
defparam sdpb_inst_3.INIT_RAM_2B = 256'h0000000000001FF8001FC0FF000000000000000000000001FCF81BFC00000000;
defparam sdpb_inst_3.INIT_RAM_2C = 256'h0000000000001FF0001FC1FF000000000000000000000000FFF81FF800000000;
defparam sdpb_inst_3.INIT_RAM_2D = 256'h0000000000001FE0001FC3DE0000000000000000000000003FF83FE000000000;
defparam sdpb_inst_3.INIT_RAM_2E = 256'h0000000000003FC0001FC3FC0000000000000000000000000FF8FF8000000000;
defparam sdpb_inst_3.INIT_RAM_2F = 256'h0000000000007FC0001FC7FC00000000000000000000000003FFFE0000000000;
defparam sdpb_inst_3.INIT_RAM_30 = 256'h000000000000FFC0001FCFF8000000000000000000000000003FE00000000000;
defparam sdpb_inst_3.INIT_RAM_31 = 256'h000000000000FFC0001FCFF00000000000000000000000000000000000000000;
defparam sdpb_inst_3.INIT_RAM_32 = 256'h000000000001FFC0001FDFE00000000000000000000000000000000000000000;
defparam sdpb_inst_3.INIT_RAM_33 = 256'h000000000003FFF0001FFFE00000000000000000000000000000000000000000;
defparam sdpb_inst_3.INIT_RAM_34 = 256'h000000000003FFFE40FFFFC00000000000000000000000000000000000000000;
defparam sdpb_inst_3.INIT_RAM_35 = 256'h000000000003FFFFFFFFFF800000000000000000000000000000000000000000;
defparam sdpb_inst_3.INIT_RAM_36 = 256'h000000000003FFFFFFFFFF000000000000000000000000000000000000000000;
defparam sdpb_inst_3.INIT_RAM_37 = 256'h000000000001FFFFFFFFFF000000000000000000000000000000000000000000;
defparam sdpb_inst_3.INIT_RAM_38 = 256'h00000000000FFF8001FFFE000000000000000000000000000000000000000000;
defparam sdpb_inst_3.INIT_RAM_39 = 256'h0000000009FFE00003FFFC000000000000000000000000000000000000000000;
defparam sdpb_inst_3.INIT_RAM_3A = 256'h00000001FFFFA803FFF0F8000000000000000000000000000000000000000000;
defparam sdpb_inst_3.INIT_RAM_3B = 256'h00000007FFFFFFFFE00000000000000000000000000000000000000000000000;
defparam sdpb_inst_3.INIT_RAM_3C = 256'h0000000011FFFFF0000000000000000000000000000000000000000000000000;
defparam sdpb_inst_3.INIT_RAM_3D = 256'h0000000000017C00000000000000000000000000000000000000000000000000;

DFFE dff_inst_0 (
  .Q(dff_q_0),
  .D(adb[14]),
  .CLK(clkb),
  .CE(ceb)
);
MUX2 mux_inst_0 (
  .O(dout[0]),
  .I0(sdpb_inst_0_dout[0]),
  .I1(sdpb_inst_1_dout[0]),
  .S0(dff_q_0)
);
MUX2 mux_inst_1 (
  .O(dout[1]),
  .I0(sdpb_inst_2_dout[1]),
  .I1(sdpb_inst_3_dout[1]),
  .S0(dff_q_0)
);
endmodule //Gowin_SDPB
